module main

fn main() {
	println('Started')
}