module argparse

pub fn new(args []string) []string {
	return
}