module video

pub fn cut_by_silence(dir string) string {
	return 'cut by silence'
}