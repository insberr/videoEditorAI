module src

fn init() {
	println('Editor initilized')
}

pub fn info() string {
	return 'Automatic video editor'
}